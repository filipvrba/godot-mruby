module src

#flag -L @VMODROOT/lib
#flag -I @VMODROOT/include/godot-headers-3.5.1
#flag -I @VMODROOT/include/mruby-3.1.0
