module src

#include <gdnative_api_struct.gen.h>
