module main

import src

fn main() {
	src.main()
}