module src

pub fn main() {

}

// [export: 'hello']
// pub fn hello() string {
//     return "Hello"
// }
