module src

pub fn main() {
	println('Hello World!')
}

[export: 'fib']
pub fn hello() string {
    return "Hello"
}
